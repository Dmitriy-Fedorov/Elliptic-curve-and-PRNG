//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Dmitriy Fedorov
// 
// Create Date:    21:25:37 11/27/2017 
// Design Name: 
// Module Name:    ROM_mod17 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
`timescale 1ns / 1ps
`define dataWidth 64
`define width 32
`define depth 32

module ROM_imod17(
	input wire[`dataWidth-1:0] readAddress,
	//input wire clk,
	output wire[`depth-1:0] data
	);
reg [`width-1:0] mem [`depth-1:0];	 //stores values for predifined modular inverse
wire [`width*2-1:0] readAddress_17;
mod17 read(
	.in(readAddress),
	.out(readAddress_17)
    );
assign data = mem[readAddress_17];
/*
always@(posedge clk)
begin
	data <= mem[readAddress];
end*/
initial
begin
	// Generated by C++ code
	mem[1] = 'd1;
	mem[2] = 'd9;
	mem[3] = 'd6;
	mem[4] = 'd13;
	mem[5] = 'd7;
	mem[6] = 'd3;
	mem[7] = 'd5;
	mem[8] = 'd15;
	mem[9] = 'd2;
	mem[10] = 'd12;
	mem[11] = 'd14;
	mem[12] = 'd10;
	mem[13] = 'd4;
	mem[14] = 'd11;
	mem[15] = 'd8;
	mem[16] = 'd16;
	
	mem[18] = 'd1;
	mem[19] = 'd9;
	mem[20] = 'd6;
	mem[21] = 'd13;
	mem[22] = 'd7;
	mem[23] = 'd3;
	mem[24] = 'd5;
	mem[25] = 'd15;
	mem[26] = 'd2;
	mem[27] = 'd12;
	mem[28] = 'd14;
	mem[29] = 'd10;
	mem[30] = 'd4;
	mem[31] = 'd11;
end
endmodule
